`ifndef __PS2_KEYBOARD_SCAN_CODES_H__
`define __PS2_KEYBOARD_SCAN_CODES_H__

`define SCANCODE_KEY_A              8'h1C
`define SCANCODE_KEY_B              8'h32
`define SCANCODE_KEY_C              8'h21
`define SCANCODE_KEY_D              8'h23
`define SCANCODE_KEY_E              8'h24
`define SCANCODE_KEY_F              8'h2B
`define SCANCODE_KEY_G              8'h34
`define SCANCODE_KEY_H              8'h33
`define SCANCODE_KEY_I              8'h43
`define SCANCODE_KEY_J              8'h3B
`define SCANCODE_KEY_K              8'h42
`define SCANCODE_KEY_L              8'h4B
`define SCANCODE_KEY_M              8'h3A
`define SCANCODE_KEY_N              8'h31
`define SCANCODE_KEY_O              8'h44
`define SCANCODE_KEY_P              8'h4D
`define SCANCODE_KEY_Q              8'h15
`define SCANCODE_KEY_R              8'h2D
`define SCANCODE_KEY_S              8'h1B
`define SCANCODE_KEY_T              8'h2C
`define SCANCODE_KEY_U              8'h3C
`define SCANCODE_KEY_V              8'h2A
`define SCANCODE_KEY_W              8'h1D
`define SCANCODE_KEY_X              8'h22
`define SCANCODE_KEY_Y              8'h35
`define SCANCODE_KEY_Z              8'h1A

`define SCANCODE_KEY_0              8'h45
`define SCANCODE_KEY_1              8'h16
`define SCANCODE_KEY_2              8'h1E
`define SCANCODE_KEY_3              8'h26
`define SCANCODE_KEY_4              8'h25
`define SCANCODE_KEY_5              8'h2E
`define SCANCODE_KEY_6              8'h36
`define SCANCODE_KEY_7              8'h3D
`define SCANCODE_KEY_8              8'h3E
`define SCANCODE_KEY_9              8'h46

`define SCANCODE_KEY_TILDE          8'h46
`define SCANCODE_KEY_MINUS          8'h4E
`define SCANCODE_KEY_EQUAL          8'h55
`define SCANCODE_KEY_BACKSLASH      8'h5D
`define SCANCODE_KEY_BACKSPACE      8'h66
`define SCANCODE_KEY_SPACE          8'h29
`define SCANCODE_KEY_TAB            8'h0D
`define SCANCODE_KEY_CAPS           8'h58

`define SCANCODE_KEY_LSHIFT         8'h12
`define SCANCODE_KEY_RSHIFT         8'h59

`define SCANCODE_KEY_LCTRL          8'h14
`define SCANCODE_KEY_LALT           8'h11

`define SCANCODE_KEY_ENTER          8'h5A
`define SCANCODE_KEY_ESCAPE         8'h76

/* --- I'm too lazy to do the F-Keys. I'll do it if the need arises. */

`endif
