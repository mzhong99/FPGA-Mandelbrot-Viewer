`ifndef __VGA_DISPLAY_H__
`define __VGA_DISPLAY_H__

`define DISP_COLS       800
`define DISP_ROWS       600
`define DISP_NPIXELS    (`DISP_COLS * `DISP_ROWS)
`define DISP_BITLEN     (`DISP_NPIXELS * 8)

`endif
